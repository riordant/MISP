LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY control_memory IS
	PORT (
		MW : OUT std_logic;
		MM : OUT std_logic;
		RW : OUT std_logic;
		MD : OUT std_logic;
		FS : OUT std_logic_vector(4 DOWNTO 0);
		MB : OUT std_logic;
		TB : OUT std_logic;
		TA : OUT std_logic;
		TD : OUT std_logic;
		PL : OUT std_logic;
		PI : OUT std_logic;
		IL : OUT std_logic;
		MC : OUT std_logic;
		MS : OUT std_logic_vector(2 DOWNTO 0);
		NA : OUT std_logic_vector(7 DOWNTO 0);
		IN_CAR : IN std_logic_vector(7 DOWNTO 0)
	);
END control_memory;
ARCHITECTURE Behavioral OF control_memory IS
	TYPE mem_array IS ARRAY(0 TO 255) OF
	std_logic_vector(27 DOWNTO 0);
BEGIN
	memory_m : PROCESS (IN_CAR)
		VARIABLE control_mem : mem_array := (
			--0
			X"000001F", -- 0 - transfer 16 0's to R0, a/b data
			outputs ALL 0'S
			X"000001F", -- 1
			X"000001F", -- 2
			X"0000000", -- 3
			X"BBBBBBB", -- 4
			X"0000000", -- 5
			X"CCCCCCC", -- 6
			X"0000000", -- 7
			X"DDDDDDD", -- 8
			X"0000000", -- 9
			X"1111111", -- A
			X"0000000", -- B
			X"2222222", -- C
			X"0000000", -- D
			X"3333333", -- E
			X"0000000", -- F
			-- 1
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 2
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 3
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 4
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 5
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 6
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 7
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 8
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- 9
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- A
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- B
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- C
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- D
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- E
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
			-- F
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000" -- F
			);
			VARIABLE addr : INTEGER;
			VARIABLE control_out : std_logic_vector(27 DOWNTO 0);
		BEGINaddr := conv_integer(IN_CAR);
			control_out := control_mem(addr);
			MW <= control_out(0);
			MM <= control_out(1);
			RW <= control_out(2);
			MD <= control_out(3);
			FS <= control_out(8 DOWNTO 4);
			MB <= control_out(9);
			TB <= control_out(10);
			TA <= control_out(11);
			TD <= control_out(12);
			PL <= control_out(13);
			PI <= control_out(14);
			IL <= control_out(15);
			MC <= control_out(16);
			MS <= control_out(19 DOWNTO 17);
			NA <= control_out(27 DOWNTO 20);
		END PROCESS;
		END Behavioral;

	