ENTITY Memory IS -- use unsigned for memory address
	PORT (
		address : IN unsigned(15 DOWNTO 0);
		write_data : IN std_logic_vector(15 DOWNTO0);
		MW : IN std_logic;
		read_data : OUT std_logic_vector(15 DOWNTO0)
	);
END Memory;
ARCHITECTURE Behavioral OF Memory IS
	TYPE mem_array IS ARRAY(0 TO 511) OF
	std_logic_vector(15 DOWNTO 0); -- define type, for
	memory arrays
BEGIN
	mem_process : PROCESS (address, write_data, MW)
		-- initialize data memory, X denotes hexadecimal number
		Variable data_mem : mem_array := (
		X"0000", X"0000", X"0003",X"0003",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000",
		X"0000", X"0000", X"0000",X"0000"
		);
		VARIABLE addr : INTEGER;
BEGIN
	addr := conv_integer(address(8 DOWNTO 0));
	IF MW = '1' THEN
		data_mem(addr) := write_data;
	ELSIF MW = '0' THEN
		read_data <= data_mem(addr) AFTER 10 ns;
	END IF;
END PROCESS;
END Behavioral;